ENTITY FULL_ADD4 IS
    PORT (
        A, B : IN BIT_VECTOR(3 DOWNTO 0);
        CIN : IN BIT;
        SUM : OUT BIT_VECTOR(3 DOWNTO 0);
        COUT : OUT BIT);
END FULL_ADD4;

ARCHITECTURE FOR_GENERATE OF FULL_ADD4 IS

    COMPONENT FULL_ADDER
        PORT (
            A, B, C : IN BIT;
            COUT, SUM : OUT BIT);
    END COMPONENT;

    SIGNAL CAR : BIT_VECTOR(4 DOWNTO 0);

BEGIN
    CAR(0) <= CIN;
    GK : FOR K IN 3 DOWNTO 0 GENERATE
        FA : FULL_ADDER PORT MAP(CAR(K), A(K), B(K), CAR(K + 1), SUM(K));
    END GENERATE GK;
    COUT <= CAR(4);
END FOR_GENERATE;