IF boolean_expression THEN
    sequential_statements
    {ELSIF boolean_expression THEN
    sequential_statements}
    [ELSE
    sequential_statements]
END IF;