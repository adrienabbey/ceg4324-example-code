FOR U0 : fa USE ENTITY work.fa(struct);