CASE expression IS
    WHEN choices => sequential_statements
    WHEN choices => sequential_statements
        [WHEN OTHERS => sequential_statements]
END CASE;