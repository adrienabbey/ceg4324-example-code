power_N := y;
WHILE i < N LOOP
    power_N := power_N * y;
END LOOP;