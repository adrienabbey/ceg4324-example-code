power_N := y;
FOR i IN 2 TO N LOOP
    power_N := power_N * y;
END LOOP;