FUNCTION identifier
    [parameter list] RETURN object TYPE IS
    subprogram declaritive items
BEGIN
    sequential statements
    RETURN expression
END [FUNCTION] identifier;