-- Chapter 2, Slide 4

ENTITY fulladder IS
    PORT (
        A, B, CIN : IN BIT;
        SUM, COUT : OUT BIT);
END fulladder;